netcdf clim_ts {
dimensions:
    xi_rho = 294 ;
    xi_u = 293 ;
    xi_v = 294 ;
    eta_rho = 194 ;
    eta_u = 194 ;
    eta_v = 193 ;
    s_rho = 32 ;
    s_w = 33 ;
    clim_time = UNLIMITED ; // (0 currently)

variables:
    float clim_time(clim_time) ;
        clim_time:long_name = "climatology clim_time" ;
        clim_time:field = "clim_time, scalar, series" ;
        clim_time:units = "days since 1940-01-01 00:00:00" ;
    float zeta(clim_time, eta_rho, xi_rho) ;
        zeta:long_name = "free-surface" ;
        zeta:units = "meter" ;
        zeta:time = "clim_time" ;
        zeta:coordinates = "lat_rho lon_rho" ;
        zeta:field = "free-surface, scalar, series" ;
    float ubar(clim_time, eta_u, xi_u) ;
        ubar:long_name = "vertically integrated u-momentum component" ;
        ubar:units = "meter second-1" ;
        ubar:time = "clim_time" ;
        ubar:coordinates = "lat_u lon_u" ;
        ubar:field = "ubar-velocity, scalar, series" ;
    float vbar(clim_time, eta_v, xi_v) ;
        vbar:long_name = "vertically integrated v-momentum component" ;
        vbar:units = "meter second-1" ;
        vbar:time = "clim_time" ;
        vbar:coordinates = "lat_v lon_v" ;
        vbar:field = "vbar-velocity, scalar, series" ;
    float u(clim_time, s_rho, eta_u, xi_u) ;
        u:long_name = "u-momentum component" ;
        u:units = "meter second-1" ;
        u:time = "clim_time" ;
        u:coordinates = "lat_u lon_u" ;
        u:field = "u-velocity, scalar, series" ;
    float v(clim_time, s_rho, eta_v, xi_v) ;
        v:long_name = "v-momentum component" ;
        v:units = "meter second-1" ;
        v:time = "clim_time" ;
        v:coordinates = "lat_v lon_v" ;
        v:field = "v-velocity, scalar, series" ;
    float temp(clim_time, s_rho, eta_rho, xi_rho) ;
        temp:long_name = "potential temperature" ;
        temp:units = "Celsius" ;
        temp:time = "clim_time" ;
        temp:coordinates = "lat_rho lon_rho" ;
        temp:field = "temperature, scalar, series" ;
    float salt(clim_time, s_rho, eta_rho, xi_rho) ;
        salt:long_name = "salinity" ;
        salt:time = "clim_time" ;
        salt:coordinates = "lat_rho lon_rho" ;
        salt:field = "salt, scalar, series" ;
    float alk(clim_time, s_rho, eta_rho, xi_rho) ;
        alk:long_name = "Alkalinity" ;
        alk:units = "mol/kg" ;
        alk:time = "clim_time" ;
        alk:coordinates = "lat_rho lon_rho" ;
        alk:field = "alk, scalar, series" ;
    float cadet_arag(clim_time, s_rho, eta_rho, xi_rho) ;
        cadet_arag:long_name = "Detrital Aragonite CaCO3" ;
        cadet_arag:units = "mol/kg" ;
        cadet_arag:time = "clim_time" ;
        cadet_arag:coordinates = "lat_rho lon_rho" ;
        cadet_arag:field = "cadet_arag, scalar, series" ;
    float cadet_calc(clim_time, s_rho, eta_rho, xi_rho) ;
        cadet_calc:long_name = "Detrital Calcite CaCO3" ;
        cadet_calc:units = "mol/kg" ;
        cadet_calc:time = "clim_time" ;
        cadet_calc:coordinates = "lat_rho lon_rho" ;
        cadet_calc:field = "cadet_calc, scalar, series" ;
    float chl(clim_time, s_rho, eta_rho, xi_rho) ;
        chl:long_name = "Chlorophyll" ;
        chl:units = "ug/kg" ;
        chl:time = "clim_time" ;
        chl:coordinates = "lat_rho lon_rho" ;
        chl:field = "dic, scalar, series" ;
    float dic(clim_time, s_rho, eta_rho, xi_rho) ;
        dic:long_name = "Dissolved Inorganic Carbon" ;
        dic:units = "mol/kg" ;
        dic:time = "clim_time" ;
        dic:coordinates = "lat_rho lon_rho" ;
        dic:field = "dic, scalar, series" ;
    float fed(clim_time, s_rho, eta_rho, xi_rho) ;
        fed:long_name = "Dissolved Iron" ;
        fed:units = "mol/kg" ;
        fed:time = "clim_time" ;
        fed:coordinates = "lat_rho lon_rho" ;
        fed:field = "fed, scalar, series" ;
    float fedet(clim_time, s_rho, eta_rho, xi_rho) ;
        fedet:long_name = "Detrital Iron" ;
        fedet:units = "mol/kg" ;
        fedet:time = "clim_time" ;
        fedet:coordinates = "lat_rho lon_rho" ;
        fedet:field = "fedet, scalar, series" ;
    float fedi(clim_time, s_rho, eta_rho, xi_rho) ;
        fedi:long_name = "Diazotroph Iron" ;
        fedi:units = "mol/kg" ;
        fedi:time = "clim_time" ;
        fedi:coordinates = "lat_rho lon_rho" ;
        fedi:field = "fedi, scalar, series" ;
    float felg(clim_time, s_rho, eta_rho, xi_rho) ;
        felg:long_name = "Large Phytoplankton Iron" ;
        felg:units = "mol/kg" ;
        felg:time = "clim_time" ;
        felg:coordinates = "lat_rho lon_rho" ;
        felg:field = "felg, scalar, series" ;
    float fesm(clim_time, s_rho, eta_rho, xi_rho) ;
        fesm:long_name = "Small Phytoplankton Iron" ;
        fesm:units = "mol/kg" ;
        fesm:time = "clim_time" ;
        fesm:coordinates = "lat_rho lon_rho" ;
        fesm:field = "fesm, scalar, series" ;
    float ldon(clim_time, s_rho, eta_rho, xi_rho) ;
        ldon:long_name = "Labile DON" ;
        ldon:units = "mol/kg" ;
        ldon:time = "clim_time" ;
        ldon:coordinates = "lat_rho lon_rho" ;
        ldon:field = "ldon, scalar, series" ;
    float ldop(clim_time, s_rho, eta_rho, xi_rho) ;
        ldop:long_name = "Labile DOP" ;
        ldop:units = "mol/kg" ;
        ldop:time = "clim_time" ;
        ldop:coordinates = "lat_rho lon_rho" ;
        ldop:field = "ldop, scalar, series" ;
    float lith(clim_time, s_rho, eta_rho, xi_rho) ;
        lith:long_name = "Lithogenic Aluminosilicate" ;
        lith:units = "g/kg" ;
        lith:time = "clim_time" ;
        lith:coordinates = "lat_rho lon_rho" ;
        lith:field = "lith, scalar, series" ;
    float lithdet(clim_time, s_rho, eta_rho, xi_rho) ;
        lithdet:long_name = "Lithogenic Aluminosilicate, detrital" ;
        lithdet:units = "g/kg" ;
        lithdet:time = "clim_time" ;
        lithdet:coordinates = "lat_rho lon_rho" ;
        lithdet:field = "lithdet, scalar, series" ;
    float nbact(clim_time, s_rho, eta_rho, xi_rho) ;
        nbact:long_name = "Bacterial Nitrogen" ;
        nbact:units = "mol/kg" ;
        nbact:time = "clim_time" ;
        nbact:coordinates = "lat_rho lon_rho" ;
        nbact:field = "nbact, scalar, series" ;
    float ndet(clim_time, s_rho, eta_rho, xi_rho) ;
        ndet:long_name = "Detrital Nitrogen" ;
        ndet:units = "mol/kg" ;
        ndet:time = "clim_time" ;
        ndet:coordinates = "lat_rho lon_rho" ;
        ndet:field = "ndet, scalar, series" ;
    float ndi(clim_time, s_rho, eta_rho, xi_rho) ;
        ndi:long_name = "Diazotroph Nitrogen" ;
        ndi:units = "mol/kg" ;
        ndi:time = "clim_time" ;
        ndi:coordinates = "lat_rho lon_rho" ;
        ndi:field = "ndi, scalar, series" ;
    float nlg(clim_time, s_rho, eta_rho, xi_rho) ;
        nlg:long_name = "Large Phytoplankton Nitrogen" ;
        nlg:units = "mol/kg" ;
        nlg:time = "clim_time" ;
        nlg:coordinates = "lat_rho lon_rho" ;
        nlg:field = "nlg, scalar, series" ;
    float nsm(clim_time, s_rho, eta_rho, xi_rho) ;
        nsm:long_name = "Small Phytoplankton Nitrogen" ;
        nsm:units = "mol/kg" ;
        nsm:time = "clim_time" ;
        nsm:coordinates = "lat_rho lon_rho" ;
        nsm:field = "nsm, scalar, series" ;
    float nh4(clim_time, s_rho, eta_rho, xi_rho) ;
        nh4:long_name = "Ammonia" ;
        nh4:units = "mol/kg" ;
        nh4:time = "clim_time" ;
        nh4:coordinates = "lat_rho lon_rho" ;
        nh4:field = "nh4, scalar, series" ;
    float no3(clim_time, s_rho, eta_rho, xi_rho) ;
        no3:long_name = "Nitrate" ;
        no3:units = "mol/kg" ;
        no3:time = "clim_time" ;
        no3:coordinates = "lat_rho lon_rho" ;
        no3:field = "no3, scalar, series" ;
    float o2(clim_time, s_rho, eta_rho, xi_rho) ;
        o2:long_name = "Oxygen" ;
        o2:units = "mol/kg" ;
        o2:time = "clim_time" ;
        o2:coordinates = "lat_rho lon_rho" ;
        o2:field = "o2, scalar, series" ;
    float pdet(clim_time, s_rho, eta_rho, xi_rho) ;
        pdet:long_name = "Detrital Phosphorus" ;
        pdet:units = "mol/kg" ;
        pdet:time = "clim_time" ;
        pdet:coordinates = "lat_rho lon_rho" ;
        pdet:field = "pdet, scalar, series" ;
    float po4(clim_time, s_rho, eta_rho, xi_rho) ;
        po4:long_name = "Phosphate" ;
        po4:units = "mol/kg" ;
        po4:time = "clim_time" ;
        po4:coordinates = "lat_rho lon_rho" ;
        po4:field = "po4, scalar, series" ;
    float srdon(clim_time, s_rho, eta_rho, xi_rho) ;
        srdon:long_name = "Semi-Refractory DON" ;
        srdon:units = "mol/kg" ;
        srdon:time = "clim_time" ;
        srdon:coordinates = "lat_rho lon_rho" ;
        srdon:field = "srdon, scalar, series" ;
    float srdop(clim_time, s_rho, eta_rho, xi_rho) ;
        srdop:long_name = "Semi-Refractory DOP" ;
        srdop:units = "mol/kg" ;
        srdop:time = "clim_time" ;
        srdop:coordinates = "lat_rho lon_rho" ;
        srdop:field = "srdop, scalar, series" ;
    float sldon(clim_time, s_rho, eta_rho, xi_rho) ;
        sldon:long_name = "Semilabile DON" ;
        sldon:units = "mol/kg" ;
        sldon:time = "clim_time" ;
        sldon:coordinates = "lat_rho lon_rho" ;
        sldon:field = "sldon, scalar, series" ;
    float sldop(clim_time, s_rho, eta_rho, xi_rho) ;
        sldop:long_name = "Semilabile DOP" ;
        sldop:units = "mol/kg" ;
        sldop:time = "clim_time" ;
        sldop:coordinates = "lat_rho lon_rho" ;
        sldop:field = "sldop, scalar, series" ;
    float sidet(clim_time, s_rho, eta_rho, xi_rho) ;
        sidet:long_name = "Detrital Silicon" ;
        sidet:units = "mol/kg" ;
        sidet:time = "clim_time" ;
        sidet:coordinates = "lat_rho lon_rho" ;
        sidet:field = "sidet, scalar, series" ;
    float silg(clim_time, s_rho, eta_rho, xi_rho) ;
        silg:long_name = "Large Phytoplankton Silicon" ;
        silg:units = "mol/kg" ;
        silg:time = "clim_time" ;
        silg:coordinates = "lat_rho lon_rho" ;
        silg:field = "silg, scalar, series" ;
    float sio4(clim_time, s_rho, eta_rho, xi_rho) ;
        sio4:long_name = "Silicate" ;
        sio4:units = "mol/kg" ;
        sio4:time = "clim_time" ;
        sio4:coordinates = "lat_rho lon_rho" ;
        sio4:field = "sio4, scalar, series" ;
    float nsmz(clim_time, s_rho, eta_rho, xi_rho) ;
        nsmz:long_name = "Small Zooplankton Nitrogen" ;
        nsmz:units = "mol/kg" ;
        nsmz:time = "clim_time" ;
        nsmz:coordinates = "lat_rho lon_rho" ;
        nsmz:field = "nsmz, scalar, series" ;
    float nmdz(clim_time, s_rho, eta_rho, xi_rho) ;
        nmdz:long_name = "Medium-sized Zooplankton Nitrogen" ;
        nmdz:units = "mol/kg" ;
        nmdz:time = "clim_time" ;
        nmdz:coordinates = "lat_rho lon_rho" ;
        nmdz:field = "nmdz, scalar, series" ;
    float nlgz(clim_time, s_rho, eta_rho, xi_rho) ;
        nlgz:long_name = "Large Zooplankton Nitrogen" ;
        nlgz:units = "mol/kg" ;
        nlgz:time = "clim_time" ;
        nlgz:coordinates = "lat_rho lon_rho" ;
        nlgz:field = "nlgz, scalar, series" ;
   float htotal(clim_time, s_rho, eta_rho, xi_rho) ;
        htotal:long_name = "H+ ion concentration" ;
        htotal:units = "mol/kg" ;
        htotal:time = "clim_time" ;
        htotal:coordinates = "lat_rho lon_rho" ;
        htotal:field = "dic, scalar, series" ;
   float irr_mem(clim_time, s_rho, eta_rho, xi_rho) ;
        irr_mem:long_name = "Irradiance memory" ;
        irr_mem:units = "Watts/m2" ;
        irr_mem:time = "clim_time" ;
        irr_mem:coordinates = "lat_rho lon_rho" ;
        irr_mem:field = "dic, scalar, series" ;
   float co3_ion(clim_time, s_rho, eta_rho, xi_rho) ;
        co3_ion:long_name = "Carbonate ion" ;
        co3_ion:units = "mol/kg" ;
        co3_ion:time = "clim_time" ;
        co3_ion:coordinates = "lat_rho lon_rho" ;
        co3_ion:field = "dic, scalar, series" ;
   float mu_mem_di(clim_time, s_rho, eta_rho, xi_rho) ;
        mu_mem_di:long_name = "Aggregation Memory Diazotrophs" ;
        mu_mem_di:units = "-" ;
        mu_mem_di:time = "clim_time" ;
        mu_mem_di:coordinates = "lat_rho lon_rho" ;
        mu_mem_di:field = "dic, scalar, series" ;
   float mu_mem_sm(clim_time, s_rho, eta_rho, xi_rho) ;
        mu_mem_sm:long_name = "Aggregation Memory Small Phyto" ;
        mu_mem_sm:units = "-" ;
        mu_mem_sm:time = "clim_time" ;
        mu_mem_sm:coordinates = "lat_rho lon_rho" ;
        mu_mem_sm:field = "dic, scalar, series" ;
   float mu_mem_lg(clim_time, s_rho, eta_rho, xi_rho) ;
        mu_mem_lg:long_name = "Aggregation Memory Large Phyto" ;
        mu_mem_lg:units = "-" ;
        mu_mem_lg:time = "clim_time" ;
        mu_mem_lg:coordinates = "lat_rho lon_rho" ;
        mu_mem_lg:field = "dic, scalar, series" ;
// global attributes:
		:title = "Climatology File" ;
		:Conventions = "CF-1.0" ;
}
