netcdf s4dvar_std_b {

dimensions:
        xi_rho = 56 ;
        eta_rho = 55 ;
        xi_u = 55 ;
        eta_u = 55 ;
        xi_v = 56 ;
        eta_v = 54 ;
        IorJ = 56 ;
        s_rho = 30 ;
        s_w = 31 ;
        boundary = 4 ;

        ocean_time = UNLIMITED ; // (0 currently)

variables:
  double ocean_time(ocean_time) ;
    ocean_time:long_name = "time since initialization" ;
    ocean_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
    ocean_time:calendar = "gregorian" ;
  double zeta_obc(ocean_time, boundary, IorJ) ;
    zeta_obc:long_name = "free-surface open boundaries standard deviation" ;
    zeta_obc:units = "meter" ;
    zeta_obc:time = "ocean_time" ;
  double ubar_obc(ocean_time, boundary, IorJ) ;
    ubar_obc:long_name = "vertically integrated u-momentum component open boundaries standard deviation" ;
    ubar_obc:units = "meter second-1" ;
    ubar_obc:time = "ocean_time" ;
  double vbar_obc(ocean_time, boundary, IorJ) ;
    vbar_obc:long_name = "vertically integrated v-momentum component open boundaries standard deviation" ;
    vbar_obc:units = "meter second-1" ;
    vbar_obc:time = "ocean_time" ;
  double u_obc(ocean_time, boundary, s_rho, IorJ) ;
    u_obc:long_name = "u-momentum component open boundaries standard deviation" ;
    u_obc:units = "meter second-1" ;
    u_obc:time = "ocean_time" ;
    u_obc:coordinates = "x_u y_u" ;
  double v_obc(ocean_time, boundary, s_rho, IorJ) ;
    v_obc:long_name = "v-momentum component open boundaries standard deviation" ;
    v_obc:units = "meter second-1" ;
    v_obc:time = "ocean_time" ;
  double temp_obc(ocean_time, boundary, s_rho, IorJ) ;
    temp_obc:long_name = "potential temperature open boundaries standard deviation" ;
    temp_obc:units = "Celsius" ;
    temp_obc:time = "ocean_time" ;
  double salt_obc(ocean_time, boundary, s_rho, IorJ) ;
    salt_obc:long_name = "salinity open boundaries standard deviation" ;
    salt_obc:time = "ocean_time" ;

// global attributes:
    :type = "ROMS/TOMS 4DVAR open boundary conditions error covariance standard deviation" ;
    :boundary_index = "West=1, South=2, East=3, North=4" ;
}
