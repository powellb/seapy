netcdf zlevel {
dimensions:
    lat = 192 ;
    lon = 382 ;
    depth = 40 ;
    time = UNLIMITED ; // (0 currently)
variables:
    float lat(lat, lon) ;
        lat:long_name = "Latitude" ;
        lat:units = "degrees_north";
    float lon(lat, lon) ;
        lon:long_name = "Longitude" ;
        lon:units = "degrees_east";
    float depth(depth) ;
        depth:long_name = "Z-Level Depth" ;
        depth:units = "meter" ;
        depth:positive = "down" ;
    float mask(lat, lon) ;
        mask:long_name = "field mask" ;
        mask:value = "0-land, 1-water" ;
    float time(time) ;
        time:long_name = "time since initialization" ;
        time:units = "hours since 1940-01-01 00:00:00" ;
    float zeta(time, lat, lon) ;
        zeta:long_name = "free-surface" ;
        zeta:units = "meter" ;
        zeta:coordinates = "lon lat" ;
        zeta:missing_value = 9.99e+10f ;
    float u(time, depth, lat, lon) ;
        u:long_name = "u-momentum component" ;
        u:units = "meter second-1" ;
        u:coordinates = "lon lat" ;
        u:missing_value = 9.99e+10f ;
    float v(time, depth, lat, lon) ;
        v:long_name = "v-momentum component" ;
        v:units = "meter second-1" ;
        v:coordinates = "lon lat" ;
        v:missing_value = 9.99e+10f ;
    float temp(time, depth, lat, lon) ;
        temp:long_name = "potential temperature" ;
        temp:units = "Celsius" ;
        temp:coordinates = "lon lat" ;
        temp:missing_value = 9.99e+10f ;
    float salt(time, depth, lat, lon) ;
        salt:long_name = "salinity" ;
        salt:units = "ppt" ;
        salt:coordinates = "lon lat" ;
        salt:missing_value = 9.99e+10f ;
// global attributes:
        :title = "Z Grid File" ;
}
