netcdf zlevel-cobalt-2d {

dimensions:
    lat = 192 ;
    lon = 382 ;
    depth = 40 ;
    time = UNLIMITED ; // (0 currently)

variables:
    float lat(lat, lon) ;
        lat:long_name = "Latitude" ;
        lat:units = "degrees_north";
    float lon(lat, lon) ;
        lon:long_name = "Longitude" ;
        lon:units = "degrees_east";
    float depth(depth) ;
        depth:long_name = "Z-Level Depth" ;
        depth:units = "meter" ;
        depth:positive = "down" ;
    float thick(depth) ;
        thick:long_name = "Z-Level Thickness" ;
        thick:units = "meter" ;
    float mask(lat, lon) ;
        mask:long_name = "field mask" ;
        mask:value = "0-land, 1-water" ;
  double time(time) ;
      time:long_name = "time since initialization" ;
      time:units = "seconds since 0000-01-01 00:00:00" ;
  float zeta(time, lat, lon) ;
      zeta:long_name = "free-surface" ;
      zeta:units = "meter" ;
      zeta:coordinates = "lon lat time" ;
  float ubar(time, lat, lon) ;
      ubar:long_name = "vertically integrated u-momentum component" ;
      ubar:units = "meter second-1" ;
      ubar:coordinates = "lon lat time" ;
  float vbar(time, lat, lon) ;
      vbar:long_name = "vertically integrated v-momentum component" ;
      vbar:units = "meter second-1" ;
      vbar:coordinates = "lon lat time" ;
  float u(time, depth, lat, lon) ;
      u:long_name = "u-momentum component" ;
      u:units = "meter second-1" ;
      u:coordinates = "lon lat depth time" ;
  float v(time, depth, lat, lon) ;
      v:long_name = "v-momentum component" ;
      v:units = "meter second-1" ;
      v:coordinates = "lon lat depth time" ;
  float temp(time, depth, lat, lon) ;
      temp:long_name = "potential temperature" ;
      temp:units = "Celsius" ;
      temp:coordinates = "lon lat depth time" ;
  float salt(time, depth, lat, lon) ;
      salt:long_name = "salinity" ;
      salt:coordinates = "lon lat depth time" ;
  float alk(time, depth, lat, lon) ;
      alk:long_name = "Alkalinity" ;
      alk:units = "mol/kg" ;
      alk:coordinates = "lon lat depth time" ;
  float cadet_arag(time, depth, lat, lon) ;
      cadet_arag:long_name = "Detrital Aragonite CaCO3" ;
      cadet_arag:units = "mol/kg" ;
      cadet_arag:coordinates = "lon lat depth time" ;
  float cadet_calc(time, depth, lat, lon) ;
      cadet_calc:long_name = "Detrital Calcite CaCO3" ;
      cadet_calc:units = "mol/kg" ;
      cadet_calc:coordinates = "lon lat depth time" ;
  float dic(time, depth, lat, lon) ;
      dic:long_name = "Dissolved Inorganic Carbon" ;
      dic:units = "mol/kg" ;
      dic:coordinates = "lon lat depth time" ;
  float fed(time, depth, lat, lon) ;
      fed:long_name = "Dissolved Iron" ;
      fed:units = "mol/kg" ;
      fed:coordinates = "lon lat depth time" ;
  float fedet(time, depth, lat, lon) ;
      fedet:long_name = "Detrital Iron" ;
      fedet:units = "mol/kg" ;
      fedet:coordinates = "lon lat depth time" ;
  float fedi(time, depth, lat, lon) ;
      fedi:long_name = "Diazotroph Iron" ;
      fedi:units = "mol/kg" ;
      fedi:coordinates = "lon lat depth time" ;
  float felg(time, depth, lat, lon) ;
      felg:long_name = "Large Phytoplankton Iron" ;
      felg:units = "mol/kg" ;
      felg:coordinates = "lon lat depth time" ;
  float fesm(time, depth, lat, lon) ;
      fesm:long_name = "Small Phytoplankton Iron" ;
      fesm:units = "mol/kg" ;
      fesm:coordinates = "lon lat depth time" ;
  float ldon(time, depth, lat, lon) ;
      ldon:long_name = "Labile DON" ;
      ldon:units = "mol/kg" ;
      ldon:coordinates = "lon lat depth time" ;
  float ldop(time, depth, lat, lon) ;
      ldop:long_name = "Labile DOP" ;
      ldop:units = "mol/kg" ;
      ldop:coordinates = "lon lat depth time" ;
  float lith(time, depth, lat, lon) ;
      lith:long_name = "Lithogenic Aluminosilicate" ;
      lith:units = "g/kg" ;
      lith:coordinates = "lon lat depth time" ;
  float lithdet(time, depth, lat, lon) ;
      lithdet:long_name = "Lithogenic Aluminosilicate, detrital" ;
      lithdet:units = "g/kg" ;
      lithdet:coordinates = "lon lat depth time" ;
  float nbact(time, depth, lat, lon) ;
      nbact:long_name = "Bacterial Nitrogen" ;
      nbact:units = "mol/kg" ;
      nbact:coordinates = "lon lat depth time" ;
  float ndet(time, depth, lat, lon) ;
      ndet:long_name = "Detrital Nitrogen" ;
      ndet:units = "mol/kg" ;
      ndet:coordinates = "lon lat depth time" ;
  float ndi(time, depth, lat, lon) ;
      ndi:long_name = "Diazotroph Nitrogen" ;
      ndi:units = "mol/kg" ;
      ndi:coordinates = "lon lat depth time" ;
  float nlg(time, depth, lat, lon) ;
      nlg:long_name = "Large Phytoplankton Nitrogen" ;
      nlg:units = "mol/kg" ;
      nlg:coordinates = "lon lat depth time" ;
  float nsm(time, depth, lat, lon) ;
      nsm:long_name = "Small Phytoplankton Nitrogen" ;
      nsm:units = "mol/kg" ;
      nsm:coordinates = "lon lat depth time" ;
  float nh4(time, depth, lat, lon) ;
      nh4:long_name = "Ammonia" ;
      nh4:units = "mol/kg" ;
      nh4:coordinates = "lon lat depth time" ;
  float no3(time, depth, lat, lon) ;
      no3:long_name = "Nitrate" ;
      no3:units = "mol/kg" ;
      no3:coordinates = "lon lat depth time" ;
  float o2(time, depth, lat, lon) ;
      o2:long_name = "Oxygen" ;
      o2:units = "mol/kg" ;
      o2:coordinates = "lon lat depth time" ;
  float pdet(time, depth, lat, lon) ;
      pdet:long_name = "Detrital Phosphorus" ;
      pdet:units = "mol/kg" ;
      pdet:coordinates = "lon lat depth time" ;
  float po4(time, depth, lat, lon) ;
      po4:long_name = "Phosphate" ;
      po4:units = "mol/kg" ;
      po4:coordinates = "lon lat depth time" ;
  float srdon(time, depth, lat, lon) ;
      srdon:long_name = "Semi-Refractory DON" ;
      srdon:units = "mol/kg" ;
      srdon:coordinates = "lon lat depth time" ;
  float srdop(time, depth, lat, lon) ;
      srdop:long_name = "Semi-Refractory DOP" ;
      srdop:units = "mol/kg" ;
      srdop:coordinates = "lon lat depth time" ;
  float sldon(time, depth, lat, lon) ;
      sldon:long_name = "Semilabile DON" ;
      sldon:units = "mol/kg" ;
      sldon:coordinates = "lon lat depth time" ;
  float sldop(time, depth, lat, lon) ;
      sldop:long_name = "Semilabile DOP" ;
      sldop:units = "mol/kg" ;
      sldop:coordinates = "lon lat depth time" ;
  float sidet(time, depth, lat, lon) ;
      sidet:long_name = "Detrital Silicon" ;
      sidet:units = "mol/kg" ;
      sidet:coordinates = "lon lat depth time" ;
  float silg(time, depth, lat, lon) ;
      silg:long_name = "Large Phytoplankton Silicon" ;
      silg:units = "mol/kg" ;
      silg:coordinates = "lon lat depth time" ;
  float sio4(time, depth, lat, lon) ;
      sio4:long_name = "Silicate" ;
      sio4:units = "mol/kg" ;
      sio4:coordinates = "lon lat depth time" ;
  float nsmz(time, depth, lat, lon) ;
      nsmz:long_name = "Small Zooplankton Nitrogen" ;
      nsmz:units = "mol/kg" ;
      nsmz:coordinates = "lon lat depth time" ;
  float nmdz(time, depth, lat, lon) ;
      nmdz:long_name = "Medium-sized Zooplankton Nitrogen" ;
      nmdz:units = "mol/kg" ;
      nmdz:coordinates = "lon lat depth time" ;
  float nlgz(time, depth, lat, lon) ;
      nlgz:long_name = "Large Zooplankton Nitrogen" ;
      nlgz:units = "mol/kg" ;
      nlgz:coordinates = "lon lat depth time" ;

// global attributes:
        :type = "Z-level output file" ;
}
