netcdf clim_ts {
dimensions:
	xi_rho = 294 ;
	xi_u = 293 ;
	xi_v = 294 ;
	eta_rho = 194 ;
	eta_u = 194 ;
	eta_v = 193 ;
	s_rho = 32 ;
	s_w = 33 ;
	clim_time = UNLIMITED ; // (0 currently)

variables:
	double clim_time(clim_time) ;
		clim_time:long_name = "climatology clim_time" ;
		clim_time:field = "clim_time, scalar, series" ;
		clim_time:units = "days since 1940-01-01 00:00:00" ;
	double zeta(clim_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:clim_time = "clim_time" ;
		zeta:coordinates = "lat_rho lon_rho" ;
		zeta:field = "free-surface, scalar, series" ;
	double ubar(clim_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:clim_time = "clim_time" ;
		ubar:coordinates = "lat_u lon_u" ;
		ubar:field = "ubar-velocity, scalar, series" ;
	double vbar(clim_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:clim_time = "clim_time" ;
		vbar:coordinates = "lat_v lon_v" ;
		vbar:field = "vbar-velocity, scalar, series" ;
	double u(clim_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:clim_time = "clim_time" ;
		u:coordinates = "lat_u lon_u" ;
		u:field = "u-velocity, scalar, series" ;
	double v(clim_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:clim_time = "clim_time" ;
		v:coordinates = "lat_v lon_v" ;
		v:field = "v-velocity, scalar, series" ;
	double temp(clim_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:clim_time = "clim_time" ;
		temp:coordinates = "lat_rho lon_rho" ;
		temp:field = "temperature, scalar, series" ;
	double salt(clim_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:clim_time = "clim_time" ;
		salt:coordinates = "lat_rho lon_rho" ;
		salt:field = "temperature, scalar, series" ;

// global attributes:
		:title = "Climatology File" ;
		:Conventions = "CF-1.0" ;
}
