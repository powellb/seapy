netcdf s4dvar_std_f {

dimensions:
        xi_rho = 56 ;
        eta_rho = 55 ;
        xi_u = 55 ;
        eta_u = 55 ;
        xi_v = 56 ;
        eta_v = 54 ;
        s_rho = 30 ;
        s_w = 31 ;
        ocean_time = UNLIMITED ; // (0 currently)

variables:
  double ocean_time(ocean_time) ;
    ocean_time:long_name = "time since initialization" ;
    ocean_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
    ocean_time:calendar = "gregorian" ;
  double sustr(ocean_time, eta_u, xi_u) ;
    sustr:long_name = "surface u-momentum stress standard deviation" ;
    sustr:units = "newton meter-2" ;
    sustr:time = "ocean_time" ;
    sustr:coordinates = "lat_u lon_u ocean_time" ;
  double svstr(ocean_time, eta_v, xi_v) ;
    svstr:long_name = "surface v-momentum stress standard deviation" ;
    svstr:units = "newton meter-2" ;
    svstr:time = "ocean_time" ;
    svstr:coordinates = "lat_v lon_v ocean_time" ;
  double shflux(ocean_time, eta_rho, xi_rho) ;
    shflux:long_name = "surface net heat flux standard deviation" ;
    shflux:units = "watt meter-2" ;
    shflux:negative_value = "upward flux, cooling" ;
    shflux:positive_value = "downward flux, heating" ;
    shflux:time = "ocean_time" ;
    shflux:coordinates = "lat_rho lon_rho ocean_time" ;
  double ssflux(ocean_time, eta_rho, xi_rho) ;
    ssflux:long_name = "surface net salt flux (E-P)*SALT standard deviation" ;
    ssflux:units = "meter second-1" ;
    ssflux:negative_value = "upward flux, freshening (net precipitation)" ;
    ssflux:positive_value = "downward flux, salting (net evaporation)" ;
    ssflux:time = "ocean_time" ;
    ssflux:coordinates = "lat_rho lon_rho ocean_time" ;

// global attributes:
    :type = "ROMS/TOMS 4DVAR surface forcing error covariance standard deviation" ;
}
