netcdf nudge_coef {
dimensions:
	xi_rho = 130 ;
	eta_rho = 82 ;
	s_rho = 36 ;
variables:
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0, 1 ;
		spherical:flag_meanings = "Cartesian spherical" ;
	float lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
		lon_rho:standard_name = "longitude" ;
	float lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
		lat_rho:standard_name = "latitude" ;
	float M2_NudgeCoef(eta_rho, xi_rho) ;
		M2_NudgeCoef:long_name = "2D momentum inverse nudging coefficients" ;
		M2_NudgeCoef:units = "day-1" ;
		M2_NudgeCoef:coordinates = "xi_rho eta_rho " ;
	float M3_NudgeCoef(s_rho, eta_rho, xi_rho) ;
		M3_NudgeCoef:long_name = "3D momentum inverse nudging coefficients" ;
		M3_NudgeCoef:units = "day-1" ;
		M3_NudgeCoef:coordinates = "xi_rho eta_rho s_rho " ;
	float temp_NudgeCoef(s_rho, eta_rho, xi_rho) ;
		temp_NudgeCoef:long_name = "temp inverse nudging coefficients" ;
		temp_NudgeCoef:units = "day-1" ;
		temp_NudgeCoef:coordinates = "xi_rho eta_rho s_rho " ;
	float salt_NudgeCoef(s_rho, eta_rho, xi_rho) ;
		salt_NudgeCoef:long_name = "salt inverse nudging coefficients" ;
		salt_NudgeCoef:units = "day-1" ;
		salt_NudgeCoef:coordinates = "xi_rho eta_rho s_rho " ;
    float alk_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        alk_NudgeCoef:long_name = "Alkalinity" ;
        alk_NudgeCoef:units = "mol/kg" ;
        alk_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float cadet_arag_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        cadet_arag_NudgeCoef:long_name = "Detrital Aragonite CaCO3" ;
        cadet_arag_NudgeCoef:units = "mol/kg" ;
        cadet_arag_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float cadet_calc_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        cadet_calc_NudgeCoef:long_name = "Detrital Calcite CaCO3" ;
        cadet_calc_NudgeCoef:units = "mol/kg" ;
        cadet_calc_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float dic_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        dic_NudgeCoef:long_name = "Dissolved Inorganic Carbon" ;
        dic_NudgeCoef:units = "mol/kg" ;
        dic_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float fed_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        fed_NudgeCoef:long_name = "Dissolved Iron" ;
        fed_NudgeCoef:units = "mol/kg" ;
        fed_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float fedet_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        fedet_NudgeCoef:long_name = "Detrital Iron" ;
        fedet_NudgeCoef:units = "mol/kg" ;
        fedet_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float fedi_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        fedi_NudgeCoef:long_name = "Diazotroph Iron" ;
        fedi_NudgeCoef:units = "mol/kg" ;
        fedi_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float felg_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        felg_NudgeCoef:long_name = "Large Phytoplankton Iron" ;
        felg_NudgeCoef:units = "mol/kg" ;
        felg_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float fesm_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        fesm_NudgeCoef:long_name = "Small Phytoplankton Iron" ;
        fesm_NudgeCoef:units = "mol/kg" ;
        fesm_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float ldon_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        ldon_NudgeCoef:long_name = "Labile DON" ;
        ldon_NudgeCoef:units = "mol/kg" ;
        ldon_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float ldop_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        ldop_NudgeCoef:long_name = "Labile DOP" ;
        ldop_NudgeCoef:units = "mol/kg" ;
        ldop_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float lith_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        lith_NudgeCoef:long_name = "Lithogenic Aluminosilicate" ;
        lith_NudgeCoef:units = "g/kg" ;
        lith_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float lithdet_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        lithdet_NudgeCoef:long_name = "Lithogenic Aluminosilicate, detrital" ;
        lithdet_NudgeCoef:units = "g/kg" ;
        lithdet_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float nbact_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        nbact_NudgeCoef:long_name = "Bacterial Nitrogen" ;
        nbact_NudgeCoef:units = "mol/kg" ;
        nbact_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float ndet_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        ndet_NudgeCoef:long_name = "Detrital Nitrogen" ;
        ndet_NudgeCoef:units = "mol/kg" ;
        ndet_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float ndi_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        ndi_NudgeCoef:long_name = "Diazotroph Nitrogen" ;
        ndi_NudgeCoef:units = "mol/kg" ;
        ndi_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float nlg_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        nlg_NudgeCoef:long_name = "Large Phytoplankton Nitrogen" ;
        nlg_NudgeCoef:units = "mol/kg" ;
        nlg_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float nsm_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        nsm_NudgeCoef:long_name = "Small Phytoplankton Nitrogen" ;
        nsm_NudgeCoef:units = "mol/kg" ;
        nsm_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float nh4_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        nh4_NudgeCoef:long_name = "Ammonia" ;
        nh4_NudgeCoef:units = "mol/kg" ;
        nh4_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float no3_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        no3_NudgeCoef:long_name = "Nitrate" ;
        no3_NudgeCoef:units = "mol/kg" ;
        no3_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float o2_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        o2_NudgeCoef:long_name = "Oxygen" ;
        o2_NudgeCoef:units = "mol/kg" ;
        o2_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float pdet_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        pdet_NudgeCoef:long_name = "Detrital Phosphorus" ;
        pdet_NudgeCoef:units = "mol/kg" ;
        pdet_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float po4_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        po4_NudgeCoef:long_name = "Phosphate" ;
        po4_NudgeCoef:units = "mol/kg" ;
        po4_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float srdon_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        srdon_NudgeCoef:long_name = "Semi-Refractory DON" ;
        srdon_NudgeCoef:units = "mol/kg" ;
        srdon_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float srdop_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        srdop_NudgeCoef:long_name = "Semi-Refractory DOP" ;
        srdop_NudgeCoef:units = "mol/kg" ;
        srdop_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float sldon_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        sldon_NudgeCoef:long_name = "Semilabile DON" ;
        sldon_NudgeCoef:units = "mol/kg" ;
        sldon_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float sldop_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        sldop_NudgeCoef:long_name = "Semilabile DOP" ;
        sldop_NudgeCoef:units = "mol/kg" ;
        sldop_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float sidet_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        sidet_NudgeCoef:long_name = "Detrital Silicon" ;
        sidet_NudgeCoef:units = "mol/kg" ;
        sidet_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float silg_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        silg_NudgeCoef:long_name = "Large Phytoplankton Silicon" ;
        silg_NudgeCoef:units = "mol/kg" ;
        silg_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float sio4_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        sio4_NudgeCoef:long_name = "Silicate" ;
        sio4_NudgeCoef:units = "mol/kg" ;
        sio4_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float nsmz_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        nsmz_NudgeCoef:long_name = "Small Zooplankton Nitrogen" ;
        nsmz_NudgeCoef:units = "mol/kg" ;
        nsmz_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float nmdz_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        nmdz_NudgeCoef:long_name = "Medium-sized Zooplankton Nitrogen" ;
        nmdz_NudgeCoef:units = "mol/kg" ;
        nmdz_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
    float nlgz_NudgeCoef(s_rho, eta_rho, xi_rho) ;
        nlgz_NudgeCoef:long_name = "Large Zooplankton Nitrogen" ;
        nlgz_NudgeCoef:units = "mol/kg" ;
        nlgz_NudgeCoef:coordinates = "lon_rho lat_rho s_rho ocean_time" ;

// global attributes:
		:type = "Nudging Coefficients file" ;
}
