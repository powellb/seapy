netcdf bry_unlimit {

dimensions:
    xi_rho = 66 ;
    eta_rho = 194 ;
    xi_u = 65 ;
    eta_u = 194 ;
    xi_v = 66 ;
    eta_v = 193 ;
    s_rho = 30 ;
    s_w = 31 ;
    bry_time = UNLIMITED ; // (0 currently)

variables:
    int spherical ;
        spherical:long_name = "grid type logical switch" ;
        spherical:flag_values = "0, 1" ;
        spherical:flag_meanings = "Cartesian spherical" ;
    int Vtransform ;
        Vtransform:long_name = "vertical terrain-following transformation equation" ;
    int Vstretching ;
        Vstretching:long_name = "vertical terrain-following stretching function" ;
    double theta_s ;
        theta_s:long_name = "S-coordinate surface control parameter" ;
    double theta_b ;
        theta_b:long_name = "S-coordinate bottom control parameter" ;
    double Tcline ;
        Tcline:long_name = "S-coordinate surface/bottom layer width" ;
        Tcline:units = "meter" ;
    double hc ;
        hc:long_name = "S-coordinate parameter, critical depth" ;
        hc:units = "meter" ;
    double s_rho(s_rho) ;
        s_rho:long_name = "S-coordinate at RHO-points" ;
        s_rho:valid_min = -1. ;
        s_rho:valid_max = 0. ;
        s_rho:positive = "up" ;
        s_rho:standard_name = "ocean_s_coordinate_g1" ;
        s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
    double s_w(s_w) ;
        s_w:long_name = "S-coordinate at W-points" ;
        s_w:valid_min = -1. ;
        s_w:valid_max = 0. ;
        s_w:positive = "up" ;
        s_w:standard_name = "ocean_s_coordinate_g1" ;
        s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
    double Cs_r(s_rho) ;
        Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
        Cs_r:valid_min = -1. ;
        Cs_r:valid_max = 0. ;
    double Cs_w(s_w) ;
        Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
        Cs_w:valid_min = -1. ;
        Cs_w:valid_max = 0. ;
    double h(eta_rho, xi_rho) ;
        h:long_name = "bathymetry at RHO-points" ;
        h:units = "meter" ;
        h:coordinates = "lon_rho lat_rho" ;
    double lon_rho(eta_rho, xi_rho) ;
        lon_rho:long_name = "longitude of RHO-points" ;
        lon_rho:units = "degree_east" ;
        lon_rho:standard_name = "longitude" ;
    double lat_rho(eta_rho, xi_rho) ;
        lat_rho:long_name = "latitude of RHO-points" ;
        lat_rho:units = "degree_north" ;
        lat_rho:standard_name = "latitude" ;
    double lon_u(eta_u, xi_u) ;
        lon_u:long_name = "longitude of U-points" ;
        lon_u:units = "degree_east" ;
        lon_u:standard_name = "longitude" ;
    double lat_u(eta_u, xi_u) ;
        lat_u:long_name = "latitude of U-points" ;
        lat_u:units = "degree_north" ;
        lat_u:standard_name = "latitude" ;
    double lon_v(eta_v, xi_v) ;
        lon_v:long_name = "longitude of V-points" ;
        lon_v:units = "degree_east" ;
        lon_v:standard_name = "longitude" ;
    double lat_v(eta_v, xi_v) ;
        lat_v:long_name = "latitude of V-points" ;
        lat_v:units = "degree_north" ;
        lat_v:standard_name = "latitude" ;
    double bry_time(bry_time) ;
        bry_time:long_name = "open boundary conditions time" ;
        bry_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
        bry_time:calendar = "gregorian" ;
    float zeta_west(bry_time, eta_rho) ;
        zeta_west:long_name = "free-surface western boundary condition" ;
        zeta_west:units = "meter" ;
        zeta_west:time = "bry_time" ;
    float zeta_east(bry_time, eta_rho) ;
        zeta_east:long_name = "free-surface eastern boundary condition" ;
        zeta_east:units = "meter" ;
        zeta_east:time = "bry_time" ;
    float zeta_south(bry_time, xi_rho) ;
        zeta_south:long_name = "free-surface southern boundary condition" ;
        zeta_south:units = "meter" ;
        zeta_south:time = "bry_time" ;
    float zeta_north(bry_time, xi_rho) ;
        zeta_north:long_name = "free-surface northern boundary condition" ;
        zeta_north:units = "meter" ;
        zeta_north:time = "bry_time" ;
    float ubar_west(bry_time, eta_u) ;
        ubar_west:long_name = "2D u-momentum western boundary condition" ;
        ubar_west:units = "meter second-1" ;
        ubar_west:time = "bry_time" ;
    float ubar_east(bry_time, eta_u) ;
        ubar_east:long_name = "2D u-momentum eastern boundary condition" ;
        ubar_east:units = "meter second-1" ;
        ubar_east:time = "bry_time" ;
    float ubar_south(bry_time, xi_u) ;
        ubar_south:long_name = "2D u-momentum southern boundary condition" ;
        ubar_south:units = "meter second-1" ;
        ubar_south:time = "bry_time" ;
    float ubar_north(bry_time, xi_u) ;
        ubar_north:long_name = "2D u-momentum northern boundary condition" ;
        ubar_north:units = "meter second-1" ;
        ubar_north:time = "bry_time" ;
    float vbar_west(bry_time, eta_v) ;
        vbar_west:long_name = "2D v-momentum western boundary condition" ;
        vbar_west:units = "meter second-1" ;
        vbar_west:time = "bry_time" ;
    float vbar_east(bry_time, eta_v) ;
        vbar_east:long_name = "2D v-momentum eastern boundary condition" ;
        vbar_east:units = "meter second-1" ;
        vbar_east:time = "bry_time" ;
    float vbar_south(bry_time, xi_v) ;
        vbar_south:long_name = "2D v-momentum southern boundary condition" ;
        vbar_south:units = "meter second-1" ;
        vbar_south:time = "bry_time" ;
    float vbar_north(bry_time, xi_v) ;
        vbar_north:long_name = "2D v-momentum northern boundary condition" ;
        vbar_north:units = "meter second-1" ;
        vbar_north:time = "bry_time" ;
    float u_west(bry_time, s_rho, eta_u) ;
        u_west:long_name = "3D u-momentum western boundary condition" ;
        u_west:units = "meter second-1" ;
        u_west:time = "bry_time" ;
    float u_east(bry_time, s_rho, eta_u) ;
        u_east:long_name = "3D u-momentum eastern boundary condition" ;
        u_east:units = "meter second-1" ;
        u_east:time = "bry_time" ;
    float u_south(bry_time, s_rho, xi_u) ;
        u_south:long_name = "3D u-momentum southern boundary condition" ;
        u_south:units = "meter second-1" ;
        u_south:time = "bry_time" ;
    float u_north(bry_time, s_rho, xi_u) ;
        u_north:long_name = "3D u-momentum northern boundary condition" ;
        u_north:units = "meter second-1" ;
        u_north:time = "bry_time" ;
    float v_west(bry_time, s_rho, eta_v) ;
        v_west:long_name = "3D v-momentum western boundary condition" ;
        v_west:units = "meter second-1" ;
        v_west:time = "bry_time" ;
    float v_east(bry_time, s_rho, eta_v) ;
        v_east:long_name = "3D v-momentum eastern boundary condition" ;
        v_east:units = "meter second-1" ;
        v_east:time = "bry_time" ;
    float v_south(bry_time, s_rho, xi_v) ;
        v_south:long_name = "3D v-momentum southern boundary condition" ;
        v_south:units = "meter second-1" ;
        v_south:time = "bry_time" ;
    float v_north(bry_time, s_rho, xi_v) ;
        v_north:long_name = "3D v-momentum northern boundary condition" ;
        v_north:units = "meter second-1" ;
        v_north:time = "bry_time" ;
    float temp_west(bry_time, s_rho, eta_rho) ;
        temp_west:long_name = "potential temperature western boundary condition" ;
        temp_west:units = "Celsius" ;
        temp_west:time = "bry_time" ;
    float temp_east(bry_time, s_rho, eta_rho) ;
        temp_east:long_name = "potential temperature eastern boundary condition" ;
        temp_east:units = "Celsius" ;
        temp_east:time = "bry_time" ;
    float temp_south(bry_time, s_rho, xi_rho) ;
        temp_south:long_name = "potential temperature southern boundary condition" ;
        temp_south:units = "Celsius" ;
        temp_south:time = "bry_time" ;
    float temp_north(bry_time, s_rho, xi_rho) ;
        temp_north:long_name = "potential temperature northern boundary condition" ;
        temp_north:units = "Celsius" ;
        temp_north:time = "bry_time" ;
    float salt_west(bry_time, s_rho, eta_rho) ;
        salt_west:long_name = "salinity western boundary condition" ;
        salt_west:time = "bry_time" ;
    float salt_east(bry_time, s_rho, eta_rho) ;
        salt_east:long_name = "salinity eastern boundary condition" ;
        salt_east:time = "bry_time" ;
    float salt_south(bry_time, s_rho, xi_rho) ;
        salt_south:long_name = "salinity southern boundary condition" ;
        salt_south:time = "bry_time" ;
    float salt_north(bry_time, s_rho, xi_rho) ;
        salt_north:long_name = "salinity northern boundary condition" ;
        salt_north:time = "bry_time" ;
    float alk_west(bry_time, s_rho, eta_rho) ;
        alk_west:long_name = "alk western boundary condition" ;
        alk_west:units = "mol/kg" ;
        alk_west:time = "bry_time" ;
    float alk_east(bry_time, s_rho, eta_rho) ;
        alk_east:long_name = "alk eastern boundary condition" ;
        alk_east:units = "mol/kg" ;
        alk_east:time = "bry_time" ;
    float alk_south(bry_time, s_rho, xi_rho) ;
        alk_south:long_name = "alk southern boundary condition" ;
        alk_south:units = "mol/kg" ;
        alk_south:time = "bry_time" ;
    float alk_north(bry_time, s_rho, xi_rho) ;
        alk_north:long_name = "alk northern boundary condition" ;
        alk_north:units = "mol/kg" ;
        alk_north:time = "bry_time" ;
    float cadet_arag_west(bry_time, s_rho, eta_rho) ;
        cadet_arag_west:long_name = "cadet_arag western boundary condition" ;
        cadet_arag_west:units = "mol/kg" ;
        cadet_arag_west:time = "bry_time" ;
    float cadet_arag_east(bry_time, s_rho, eta_rho) ;
        cadet_arag_east:long_name = "cadet_arag eastern boundary condition" ;
        cadet_arag_east:units = "mol/kg" ;
        cadet_arag_east:time = "bry_time" ;
    float cadet_arag_south(bry_time, s_rho, xi_rho) ;
        cadet_arag_south:long_name = "cadet_arag southern boundary condition" ;
        cadet_arag_south:units = "mol/kg" ;
        cadet_arag_south:time = "bry_time" ;
    float cadet_arag_north(bry_time, s_rho, xi_rho) ;
        cadet_arag_north:long_name = "cadet_arag northern boundary condition" ;
        cadet_arag_north:units = "mol/kg" ;
        cadet_arag_north:time = "bry_time" ;
    float cadet_calc_west(bry_time, s_rho, eta_rho) ;
        cadet_calc_west:long_name = "cadet_calc western boundary condition" ;
        cadet_calc_west:units = "mol/kg" ;
        cadet_calc_west:time = "bry_time" ;
    float cadet_calc_east(bry_time, s_rho, eta_rho) ;
        cadet_calc_east:long_name = "cadet_calc eastern boundary condition" ;
        cadet_calc_east:units = "mol/kg" ;
        cadet_calc_east:time = "bry_time" ;
    float cadet_calc_south(bry_time, s_rho, xi_rho) ;
        cadet_calc_south:long_name = "cadet_calc southern boundary condition" ;
        cadet_calc_south:units = "mol/kg" ;
        cadet_calc_south:time = "bry_time" ;
    float cadet_calc_north(bry_time, s_rho, xi_rho) ;
        cadet_calc_north:long_name = "cadet_calc northern boundary condition" ;
        cadet_calc_north:units = "mol/kg" ;
        cadet_calc_north:time = "bry_time" ;
    float dic_west(bry_time, s_rho, eta_rho) ;
        dic_west:long_name = "dic western boundary condition" ;
        dic_west:units = "mol/kg" ;
        dic_west:time = "bry_time" ;
    float dic_east(bry_time, s_rho, eta_rho) ;
        dic_east:long_name = "dic eastern boundary condition" ;
        dic_east:units = "mol/kg" ;
        dic_east:time = "bry_time" ;
    float dic_south(bry_time, s_rho, xi_rho) ;
        dic_south:long_name = "dic southern boundary condition" ;
        dic_south:units = "mol/kg" ;
        dic_south:time = "bry_time" ;
    float dic_north(bry_time, s_rho, xi_rho) ;
        dic_north:long_name = "dic northern boundary condition" ;
        dic_north:units = "mol/kg" ;
        dic_north:time = "bry_time" ;
    float fed_west(bry_time, s_rho, eta_rho) ;
        fed_west:long_name = "fed western boundary condition" ;
        fed_west:units = "mol/kg" ;
        fed_west:time = "bry_time" ;
    float fed_east(bry_time, s_rho, eta_rho) ;
        fed_east:long_name = "fed eastern boundary condition" ;
        fed_east:units = "mol/kg" ;
        fed_east:time = "bry_time" ;
    float fed_south(bry_time, s_rho, xi_rho) ;
        fed_south:long_name = "fed southern boundary condition" ;
        fed_south:units = "mol/kg" ;
        fed_south:time = "bry_time" ;
    float fed_north(bry_time, s_rho, xi_rho) ;
        fed_north:long_name = "fed northern boundary condition" ;
        fed_north:units = "mol/kg" ;
        fed_north:time = "bry_time" ;
    float fedet_west(bry_time, s_rho, eta_rho) ;
        fedet_west:long_name = "fedet western boundary condition" ;
        fedet_west:units = "mol/kg" ;
        fedet_west:time = "bry_time" ;
    float fedet_east(bry_time, s_rho, eta_rho) ;
        fedet_east:long_name = "fedet eastern boundary condition" ;
        fedet_east:units = "mol/kg" ;
        fedet_east:time = "bry_time" ;
    float fedet_south(bry_time, s_rho, xi_rho) ;
        fedet_south:long_name = "fedet southern boundary condition" ;
        fedet_south:units = "mol/kg" ;
        fedet_south:time = "bry_time" ;
    float fedet_north(bry_time, s_rho, xi_rho) ;
        fedet_north:long_name = "fedet northern boundary condition" ;
        fedet_north:units = "mol/kg" ;
        fedet_north:time = "bry_time" ;
    float fedi_west(bry_time, s_rho, eta_rho) ;
        fedi_west:long_name = "fedi western boundary condition" ;
        fedi_west:units = "mol/kg" ;
        fedi_west:time = "bry_time" ;
    float fedi_east(bry_time, s_rho, eta_rho) ;
        fedi_east:long_name = "fedi eastern boundary condition" ;
        fedi_east:units = "mol/kg" ;
        fedi_east:time = "bry_time" ;
    float fedi_south(bry_time, s_rho, xi_rho) ;
        fedi_south:long_name = "fedi southern boundary condition" ;
        fedi_south:units = "mol/kg" ;
        fedi_south:time = "bry_time" ;
    float fedi_north(bry_time, s_rho, xi_rho) ;
        fedi_north:long_name = "fedi northern boundary condition" ;
        fedi_north:units = "mol/kg" ;
        fedi_north:time = "bry_time" ;
    float felg_west(bry_time, s_rho, eta_rho) ;
        felg_west:long_name = "felg western boundary condition" ;
        felg_west:units = "mol/kg" ;
        felg_west:time = "bry_time" ;
    float felg_east(bry_time, s_rho, eta_rho) ;
        felg_east:long_name = "felg eastern boundary condition" ;
        felg_east:units = "mol/kg" ;
        felg_east:time = "bry_time" ;
    float felg_south(bry_time, s_rho, xi_rho) ;
        felg_south:long_name = "felg southern boundary condition" ;
        felg_south:units = "mol/kg" ;
        felg_south:time = "bry_time" ;
    float felg_north(bry_time, s_rho, xi_rho) ;
        felg_north:long_name = "felg northern boundary condition" ;
        felg_north:units = "mol/kg" ;
        felg_north:time = "bry_time" ;
    float fesm_west(bry_time, s_rho, eta_rho) ;
        fesm_west:long_name = "fesm western boundary condition" ;
        fesm_west:units = "mol/kg" ;
        fesm_west:time = "bry_time" ;
    float fesm_east(bry_time, s_rho, eta_rho) ;
        fesm_east:long_name = "fesm eastern boundary condition" ;
        fesm_east:units = "mol/kg" ;
        fesm_east:time = "bry_time" ;
    float fesm_south(bry_time, s_rho, xi_rho) ;
        fesm_south:long_name = "fesm southern boundary condition" ;
        fesm_south:units = "mol/kg" ;
        fesm_south:time = "bry_time" ;
    float fesm_north(bry_time, s_rho, xi_rho) ;
        fesm_north:long_name = "fesm northern boundary condition" ;
        fesm_north:units = "mol/kg" ;
        fesm_north:time = "bry_time" ;
    float ldon_west(bry_time, s_rho, eta_rho) ;
        ldon_west:long_name = "ldon western boundary condition" ;
        ldon_west:units = "mol/kg" ;
        ldon_west:time = "bry_time" ;
    float ldon_east(bry_time, s_rho, eta_rho) ;
        ldon_east:long_name = "ldon eastern boundary condition" ;
        ldon_east:units = "mol/kg" ;
        ldon_east:time = "bry_time" ;
    float ldon_south(bry_time, s_rho, xi_rho) ;
        ldon_south:long_name = "ldon southern boundary condition" ;
        ldon_south:units = "mol/kg" ;
        ldon_south:time = "bry_time" ;
    float ldon_north(bry_time, s_rho, xi_rho) ;
        ldon_north:long_name = "ldon northern boundary condition" ;
        ldon_north:units = "mol/kg" ;
        ldon_north:time = "bry_time" ;
    float ldop_west(bry_time, s_rho, eta_rho) ;
        ldop_west:long_name = "ldop western boundary condition" ;
        ldop_west:units = "mol/kg" ;
        ldop_west:time = "bry_time" ;
    float ldop_east(bry_time, s_rho, eta_rho) ;
        ldop_east:long_name = "ldop eastern boundary condition" ;
        ldop_east:units = "mol/kg" ;
        ldop_east:time = "bry_time" ;
    float ldop_south(bry_time, s_rho, xi_rho) ;
        ldop_south:long_name = "ldop southern boundary condition" ;
        ldop_south:units = "mol/kg" ;
        ldop_south:time = "bry_time" ;
    float ldop_north(bry_time, s_rho, xi_rho) ;
        ldop_north:long_name = "ldop northern boundary condition" ;
        ldop_north:units = "mol/kg" ;
        ldop_north:time = "bry_time" ;
    float lith_west(bry_time, s_rho, eta_rho) ;
        lith_west:long_name = "lith western boundary condition" ;
        lith_west:units = "g/kg" ;
        lith_west:time = "bry_time" ;
    float lith_east(bry_time, s_rho, eta_rho) ;
        lith_east:long_name = "lith eastern boundary condition" ;
        lith_east:units = "g/kg" ;
        lith_east:time = "bry_time" ;
    float lith_south(bry_time, s_rho, xi_rho) ;
        lith_south:long_name = "lith southern boundary condition" ;
        lith_south:units = "g/kg" ;
        lith_south:time = "bry_time" ;
    float lith_north(bry_time, s_rho, xi_rho) ;
        lith_north:long_name = "lith northern boundary condition" ;
        lith_north:units = "g/kg" ;
        lith_north:time = "bry_time" ;
    float lithdet_west(bry_time, s_rho, eta_rho) ;
        lithdet_west:long_name = "lithdet western boundary condition" ;
        lithdet_west:units = "g/kg" ;
        lithdet_west:time = "bry_time" ;
    float lithdet_east(bry_time, s_rho, eta_rho) ;
        lithdet_east:long_name = "lithdet eastern boundary condition" ;
        lithdet_east:units = "g/kg" ;
        lithdet_east:time = "bry_time" ;
    float lithdet_south(bry_time, s_rho, xi_rho) ;
        lithdet_south:long_name = "lithdet southern boundary condition" ;
        lithdet_south:units = "g/kg" ;
        lithdet_south:time = "bry_time" ;
    float lithdet_north(bry_time, s_rho, xi_rho) ;
        lithdet_north:long_name = "lithdet northern boundary condition" ;
        lithdet_north:units = "g/kg" ;
        lithdet_north:time = "bry_time" ;
    float nbact_west(bry_time, s_rho, eta_rho) ;
        nbact_west:long_name = "nbact western boundary condition" ;
        nbact_west:units = "mol/kg" ;
        nbact_west:time = "bry_time" ;
    float nbact_east(bry_time, s_rho, eta_rho) ;
        nbact_east:long_name = "nbact eastern boundary condition" ;
        nbact_east:units = "mol/kg" ;
        nbact_east:time = "bry_time" ;
    float nbact_south(bry_time, s_rho, xi_rho) ;
        nbact_south:long_name = "nbact southern boundary condition" ;
        nbact_south:units = "mol/kg" ;
        nbact_south:time = "bry_time" ;
    float nbact_north(bry_time, s_rho, xi_rho) ;
        nbact_north:long_name = "nbact northern boundary condition" ;
        nbact_north:units = "mol/kg" ;
        nbact_north:time = "bry_time" ;
    float ndet_west(bry_time, s_rho, eta_rho) ;
        ndet_west:long_name = "ndet western boundary condition" ;
        ndet_west:units = "mol/kg" ;
        ndet_west:time = "bry_time" ;
    float ndet_east(bry_time, s_rho, eta_rho) ;
        ndet_east:long_name = "ndet eastern boundary condition" ;
        ndet_east:units = "mol/kg" ;
        ndet_east:time = "bry_time" ;
    float ndet_south(bry_time, s_rho, xi_rho) ;
        ndet_south:long_name = "ndet southern boundary condition" ;
        ndet_south:units = "mol/kg" ;
        ndet_south:time = "bry_time" ;
    float ndet_north(bry_time, s_rho, xi_rho) ;
        ndet_north:long_name = "ndet northern boundary condition" ;
        ndet_north:units = "mol/kg" ;
        ndet_north:time = "bry_time" ;
    float ndi_west(bry_time, s_rho, eta_rho) ;
        ndi_west:long_name = "ndi western boundary condition" ;
        ndi_west:units = "mol/kg" ;
        ndi_west:time = "bry_time" ;
    float ndi_east(bry_time, s_rho, eta_rho) ;
        ndi_east:long_name = "ndi eastern boundary condition" ;
        ndi_east:units = "mol/kg" ;
        ndi_east:time = "bry_time" ;
    float ndi_south(bry_time, s_rho, xi_rho) ;
        ndi_south:long_name = "ndi southern boundary condition" ;
        ndi_south:units = "mol/kg" ;
        ndi_south:time = "bry_time" ;
    float ndi_north(bry_time, s_rho, xi_rho) ;
        ndi_north:long_name = "ndi northern boundary condition" ;
        ndi_north:units = "mol/kg" ;
        ndi_north:time = "bry_time" ;
    float nlg_west(bry_time, s_rho, eta_rho) ;
        nlg_west:long_name = "nlg western boundary condition" ;
        nlg_west:units = "mol/kg" ;
        nlg_west:time = "bry_time" ;
    float nlg_east(bry_time, s_rho, eta_rho) ;
        nlg_east:long_name = "nlg eastern boundary condition" ;
        nlg_east:units = "mol/kg" ;
        nlg_east:time = "bry_time" ;
    float nlg_south(bry_time, s_rho, xi_rho) ;
        nlg_south:long_name = "nlg southern boundary condition" ;
        nlg_south:units = "mol/kg" ;
        nlg_south:time = "bry_time" ;
    float nlg_north(bry_time, s_rho, xi_rho) ;
        nlg_north:long_name = "nlg northern boundary condition" ;
        nlg_north:units = "mol/kg" ;
        nlg_north:time = "bry_time" ;
    float nsm_west(bry_time, s_rho, eta_rho) ;
        nsm_west:long_name = "nsm western boundary condition" ;
        nsm_west:units = "mol/kg" ;
        nsm_west:time = "bry_time" ;
    float nsm_east(bry_time, s_rho, eta_rho) ;
        nsm_east:long_name = "nsm eastern boundary condition" ;
        nsm_east:units = "mol/kg" ;
        nsm_east:time = "bry_time" ;
    float nsm_south(bry_time, s_rho, xi_rho) ;
        nsm_south:long_name = "nsm southern boundary condition" ;
        nsm_south:units = "mol/kg" ;
        nsm_south:time = "bry_time" ;
    float nsm_north(bry_time, s_rho, xi_rho) ;
        nsm_north:long_name = "nsm northern boundary condition" ;
        nsm_north:units = "mol/kg" ;
        nsm_north:time = "bry_time" ;
    float nh4_west(bry_time, s_rho, eta_rho) ;
        nh4_west:long_name = "nh4 western boundary condition" ;
        nh4_west:units = "mol/kg" ;
        nh4_west:time = "bry_time" ;
    float nh4_east(bry_time, s_rho, eta_rho) ;
        nh4_east:long_name = "nh4 eastern boundary condition" ;
        nh4_east:units = "mol/kg" ;
        nh4_east:time = "bry_time" ;
    float nh4_south(bry_time, s_rho, xi_rho) ;
        nh4_south:long_name = "nh4 southern boundary condition" ;
        nh4_south:units = "mol/kg" ;
        nh4_south:time = "bry_time" ;
    float nh4_north(bry_time, s_rho, xi_rho) ;
        nh4_north:long_name = "nh4 northern boundary condition" ;
        nh4_north:units = "mol/kg" ;
        nh4_north:time = "bry_time" ;
    float no3_west(bry_time, s_rho, eta_rho) ;
        no3_west:long_name = "no3 western boundary condition" ;
        no3_west:units = "mol/kg" ;
        no3_west:time = "bry_time" ;
    float no3_east(bry_time, s_rho, eta_rho) ;
        no3_east:long_name = "no3 eastern boundary condition" ;
        no3_east:units = "mol/kg" ;
        no3_east:time = "bry_time" ;
    float no3_south(bry_time, s_rho, xi_rho) ;
        no3_south:long_name = "no3 southern boundary condition" ;
        no3_south:units = "mol/kg" ;
        no3_south:time = "bry_time" ;
    float no3_north(bry_time, s_rho, xi_rho) ;
        no3_north:long_name = "no3 northern boundary condition" ;
        no3_north:units = "mol/kg" ;
        no3_north:time = "bry_time" ;
    float o2_west(bry_time, s_rho, eta_rho) ;
        o2_west:long_name = "o2 western boundary condition" ;
        o2_west:units = "mol/kg" ;
        o2_west:time = "bry_time" ;
    float o2_east(bry_time, s_rho, eta_rho) ;
        o2_east:long_name = "o2 eastern boundary condition" ;
        o2_east:units = "mol/kg" ;
        o2_east:time = "bry_time" ;
    float o2_south(bry_time, s_rho, xi_rho) ;
        o2_south:long_name = "o2 southern boundary condition" ;
        o2_south:units = "mol/kg" ;
        o2_south:time = "bry_time" ;
    float o2_north(bry_time, s_rho, xi_rho) ;
        o2_north:long_name = "o2 northern boundary condition" ;
        o2_north:units = "mol/kg" ;
        o2_north:time = "bry_time" ;
    float pdet_west(bry_time, s_rho, eta_rho) ;
        pdet_west:long_name = "pdet western boundary condition" ;
        pdet_west:units = "mol/kg" ;
        pdet_west:time = "bry_time" ;
    float pdet_east(bry_time, s_rho, eta_rho) ;
        pdet_east:long_name = "pdet eastern boundary condition" ;
        pdet_east:units = "mol/kg" ;
        pdet_east:time = "bry_time" ;
    float pdet_south(bry_time, s_rho, xi_rho) ;
        pdet_south:long_name = "pdet southern boundary condition" ;
        pdet_south:units = "mol/kg" ;
        pdet_south:time = "bry_time" ;
    float pdet_north(bry_time, s_rho, xi_rho) ;
        pdet_north:long_name = "pdet northern boundary condition" ;
        pdet_north:units = "mol/kg" ;
        pdet_north:time = "bry_time" ;
    float po4_west(bry_time, s_rho, eta_rho) ;
        po4_west:long_name = "po4 western boundary condition" ;
        po4_west:units = "mol/kg" ;
        po4_west:time = "bry_time" ;
    float po4_east(bry_time, s_rho, eta_rho) ;
        po4_east:long_name = "po4 eastern boundary condition" ;
        po4_east:units = "mol/kg" ;
        po4_east:time = "bry_time" ;
    float po4_south(bry_time, s_rho, xi_rho) ;
        po4_south:long_name = "po4 southern boundary condition" ;
        po4_south:units = "mol/kg" ;
        po4_south:time = "bry_time" ;
    float po4_north(bry_time, s_rho, xi_rho) ;
        po4_north:long_name = "po4 northern boundary condition" ;
        po4_north:units = "mol/kg" ;
        po4_north:time = "bry_time" ;
    float srdon_west(bry_time, s_rho, eta_rho) ;
        srdon_west:long_name = "srdon western boundary condition" ;
        srdon_west:units = "mol/kg" ;
        srdon_west:time = "bry_time" ;
    float srdon_east(bry_time, s_rho, eta_rho) ;
        srdon_east:long_name = "srdon eastern boundary condition" ;
        srdon_east:units = "mol/kg" ;
        srdon_east:time = "bry_time" ;
    float srdon_south(bry_time, s_rho, xi_rho) ;
        srdon_south:long_name = "srdon southern boundary condition" ;
        srdon_south:units = "mol/kg" ;
        srdon_south:time = "bry_time" ;
    float srdon_north(bry_time, s_rho, xi_rho) ;
        srdon_north:long_name = "srdon northern boundary condition" ;
        srdon_north:units = "mol/kg" ;
        srdon_north:time = "bry_time" ;
    float srdop_west(bry_time, s_rho, eta_rho) ;
        srdop_west:long_name = "srdop western boundary condition" ;
        srdop_west:units = "mol/kg" ;
        srdop_west:time = "bry_time" ;
    float srdop_east(bry_time, s_rho, eta_rho) ;
        srdop_east:long_name = "srdop eastern boundary condition" ;
        srdop_east:units = "mol/kg" ;
        srdop_east:time = "bry_time" ;
    float srdop_south(bry_time, s_rho, xi_rho) ;
        srdop_south:long_name = "srdop southern boundary condition" ;
        srdop_south:units = "mol/kg" ;
        srdop_south:time = "bry_time" ;
    float srdop_north(bry_time, s_rho, xi_rho) ;
        srdop_north:long_name = "srdop northern boundary condition" ;
        srdop_north:units = "mol/kg" ;
        srdop_north:time = "bry_time" ;
    float sldon_west(bry_time, s_rho, eta_rho) ;
        sldon_west:long_name = "sldon western boundary condition" ;
        sldon_west:units = "mol/kg" ;
        sldon_west:time = "bry_time" ;
    float sldon_east(bry_time, s_rho, eta_rho) ;
        sldon_east:long_name = "sldon eastern boundary condition" ;
        sldon_east:units = "mol/kg" ;
        sldon_east:time = "bry_time" ;
    float sldon_south(bry_time, s_rho, xi_rho) ;
        sldon_south:long_name = "sldon southern boundary condition" ;
        sldon_south:units = "mol/kg" ;
        sldon_south:time = "bry_time" ;
    float sldon_north(bry_time, s_rho, xi_rho) ;
        sldon_north:long_name = "sldon northern boundary condition" ;
        sldon_north:units = "mol/kg" ;
        sldon_north:time = "bry_time" ;
    float sldop_west(bry_time, s_rho, eta_rho) ;
        sldop_west:long_name = "sldop western boundary condition" ;
        sldop_west:units = "mol/kg" ;
        sldop_west:time = "bry_time" ;
    float sldop_east(bry_time, s_rho, eta_rho) ;
        sldop_east:long_name = "sldop eastern boundary condition" ;
        sldop_east:units = "mol/kg" ;
        sldop_east:time = "bry_time" ;
    float sldop_south(bry_time, s_rho, xi_rho) ;
        sldop_south:long_name = "sldop southern boundary condition" ;
        sldop_south:units = "mol/kg" ;
        sldop_south:time = "bry_time" ;
    float sldop_north(bry_time, s_rho, xi_rho) ;
        sldop_north:long_name = "sldop northern boundary condition" ;
        sldop_north:units = "mol/kg" ;
        sldop_north:time = "bry_time" ;
    float sidet_west(bry_time, s_rho, eta_rho) ;
        sidet_west:long_name = "sidet western boundary condition" ;
        sidet_west:units = "mol/kg" ;
        sidet_west:time = "bry_time" ;
    float sidet_east(bry_time, s_rho, eta_rho) ;
        sidet_east:long_name = "sidet eastern boundary condition" ;
        sidet_east:units = "mol/kg" ;
        sidet_east:time = "bry_time" ;
    float sidet_south(bry_time, s_rho, xi_rho) ;
        sidet_south:long_name = "sidet southern boundary condition" ;
        sidet_south:units = "mol/kg" ;
        sidet_south:time = "bry_time" ;
    float sidet_north(bry_time, s_rho, xi_rho) ;
        sidet_north:long_name = "sidet northern boundary condition" ;
        sidet_north:units = "mol/kg" ;
        sidet_north:time = "bry_time" ;
    float silg_west(bry_time, s_rho, eta_rho) ;
        silg_west:long_name = "silg western boundary condition" ;
        silg_west:units = "mol/kg" ;
        silg_west:time = "bry_time" ;
    float silg_east(bry_time, s_rho, eta_rho) ;
        silg_east:long_name = "silg eastern boundary condition" ;
        silg_east:units = "mol/kg" ;
        silg_east:time = "bry_time" ;
    float silg_south(bry_time, s_rho, xi_rho) ;
        silg_south:long_name = "silg southern boundary condition" ;
        silg_south:units = "mol/kg" ;
        silg_south:time = "bry_time" ;
    float silg_north(bry_time, s_rho, xi_rho) ;
        silg_north:long_name = "silg northern boundary condition" ;
        silg_north:units = "mol/kg" ;
        silg_north:time = "bry_time" ;
    float sio4_west(bry_time, s_rho, eta_rho) ;
        sio4_west:long_name = "sio4 western boundary condition" ;
        sio4_west:units = "mol/kg" ;
        sio4_west:time = "bry_time" ;
    float sio4_east(bry_time, s_rho, eta_rho) ;
        sio4_east:long_name = "sio4 eastern boundary condition" ;
        sio4_east:units = "mol/kg" ;
        sio4_east:time = "bry_time" ;
    float sio4_south(bry_time, s_rho, xi_rho) ;
        sio4_south:long_name = "sio4 southern boundary condition" ;
        sio4_south:units = "mol/kg" ;
        sio4_south:time = "bry_time" ;
    float sio4_north(bry_time, s_rho, xi_rho) ;
        sio4_north:long_name = "sio4 northern boundary condition" ;
        sio4_north:units = "mol/kg" ;
        sio4_north:time = "bry_time" ;
    float nsmz_west(bry_time, s_rho, eta_rho) ;
        nsmz_west:long_name = "nsmz western boundary condition" ;
        nsmz_west:units = "mol/kg" ;
        nsmz_west:time = "bry_time" ;
    float nsmz_east(bry_time, s_rho, eta_rho) ;
        nsmz_east:long_name = "nsmz eastern boundary condition" ;
        nsmz_east:units = "mol/kg" ;
        nsmz_east:time = "bry_time" ;
    float nsmz_south(bry_time, s_rho, xi_rho) ;
        nsmz_south:long_name = "nsmz southern boundary condition" ;
        nsmz_south:units = "mol/kg" ;
        nsmz_south:time = "bry_time" ;
    float nsmz_north(bry_time, s_rho, xi_rho) ;
        nsmz_north:long_name = "nsmz northern boundary condition" ;
        nsmz_north:units = "mol/kg" ;
        nsmz_north:time = "bry_time" ;
    float nmdz_west(bry_time, s_rho, eta_rho) ;
        nmdz_west:long_name = "nmdz western boundary condition" ;
        nmdz_west:units = "mol/kg" ;
        nmdz_west:time = "bry_time" ;
    float nmdz_east(bry_time, s_rho, eta_rho) ;
        nmdz_east:long_name = "nmdz eastern boundary condition" ;
        nmdz_east:units = "mol/kg" ;
        nmdz_east:time = "bry_time" ;
    float nmdz_south(bry_time, s_rho, xi_rho) ;
        nmdz_south:long_name = "nmdz southern boundary condition" ;
        nmdz_south:units = "mol/kg" ;
        nmdz_south:time = "bry_time" ;
    float nmdz_north(bry_time, s_rho, xi_rho) ;
        nmdz_north:long_name = "nmdz northern boundary condition" ;
        nmdz_north:units = "mol/kg" ;
        nmdz_north:time = "bry_time" ;
    float nlgz_west(bry_time, s_rho, eta_rho) ;
        nlgz_west:long_name = "nlgz western boundary condition" ;
        nlgz_west:units = "mol/kg" ;
        nlgz_west:time = "bry_time" ;
    float nlgz_east(bry_time, s_rho, eta_rho) ;
        nlgz_east:long_name = "nlgz eastern boundary condition" ;
        nlgz_east:units = "mol/kg" ;
        nlgz_east:time = "bry_time" ;
    float nlgz_south(bry_time, s_rho, xi_rho) ;
        nlgz_south:long_name = "nlgz southern boundary condition" ;
        nlgz_south:units = "mol/kg" ;
        nlgz_south:time = "bry_time" ;
    float nlgz_north(bry_time, s_rho, xi_rho) ;
        nlgz_north:long_name = "nlgz northern boundary condition" ;
        nlgz_north:units = "mol/kg" ;
        nlgz_north:time = "bry_time" ;
// global attributes:
		:type = "BOUNDARY FORCING" ;
}
