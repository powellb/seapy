netcdf roms_grid {
dimensions:
	xi_psi = 293 ;
	xi_rho = 294 ;
	xi_u = 293 ;
	xi_v = 294 ;
	eta_psi = 193 ;
	eta_rho = 194 ;
	eta_u = 194 ;
	eta_v = 193 ;
	two = 2 ;

variables:
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	char JPRJ(two) ;
		JPRJ:long_name = "Map projection type" ;
		JPRJ:option\(ME\) = "Mercator" ;
		JPRJ:option\(ST\) = "Stereographic" ;
		JPRJ:option\(LC\) = "Lambert conformal conic" ;
	float PLAT(two) ;
		PLAT:long_name = "Reference latitude(s) for map projection" ;
		PLAT:units = "degree_north" ;
	float PLONG ;
		PLONG:long_name = "Reference longitude for map projection" ;
		PLONG:units = "degree_east" ;
	float ROTA ;
		ROTA:long_name = "Rotation angle for map projection" ;
		ROTA:units = "degree" ;
	char JLTS(two) ;
		JLTS:long_name = "How limits of map are chosen" ;
		JLTS:option\(CO\) = "P1, .. P4 define two opposite corners " ;
		JLTS:option\(MA\) = "Maximum (whole world)" ;
		JLTS:option\(AN\) = "Angles - P1..P4 define angles to edge of domain" ;
		JLTS:option\(LI\) = "Limits - P1..P4 define limits in u,v space" ;
	float P1 ;
		P1:long_name = "Map limit parameter number 1" ;
	float P2 ;
		P2:long_name = "Map limit parameter number 2" ;
	float P3 ;
		P3:long_name = "Map limit parameter number 3" ;
	float P4 ;
		P4:long_name = "Map limit parameter number 4" ;
	float XOFF ;
		XOFF:long_name = "Offset in x direction" ;
		XOFF:units = "meter" ;
	float YOFF ;
		YOFF:long_name = "Offset in y direction" ;
		YOFF:units = "meter" ;
	short depthmin ;
		depthmin:long_name = "Shallow bathymetry clipping depth" ;
		depthmin:units = "meter" ;
	short depthmax ;
		depthmax:long_name = "Deep bathymetry clipping depth" ;
		depthmax:units = "meter" ;
	char spherical ;
		spherical:long_name = "Grid type logical switch" ;
		spherical:option\(T\) = "spherical" ;
		spherical:option\(F\) = "Cartesian" ;
	double hraw(eta_rho, xi_rho) ;
		hraw:long_name = "Working bathymetry at RHO-points" ;
		hraw:units = "meter" ;
		hraw:field = "bath, scalar" ;
	double h(eta_rho, xi_rho) ;
		h:long_name = "Final bathymetry at RHO-points" ;
		h:units = "meter" ;
		h:field = "bath, scalar" ;
	double f(eta_rho, xi_rho) ;
		f:long_name = "Coriolis parameter at RHO-points" ;
		f:units = "second-1" ;
		f:field = "Coriolis, scalar" ;
	double pm(eta_rho, xi_rho) ;
		pm:long_name = "curvilinear coordinate metric in XI" ;
		pm:units = "meter-1" ;
		pm:field = "pm, scalar" ;
	double pn(eta_rho, xi_rho) ;
		pn:long_name = "curvilinear coordinate metric in ETA" ;
		pn:units = "meter-1" ;
		pn:field = "pn, scalar" ;
	double dndx(eta_rho, xi_rho) ;
		dndx:long_name = "xi derivative of inverse metric factor pn" ;
		dndx:units = "meter" ;
		dndx:field = "dndx, scalar" ;
	double dmde(eta_rho, xi_rho) ;
		dmde:long_name = "eta derivative of inverse metric factor pm" ;
		dmde:units = "meter" ;
		dmde:field = "dmde, scalar" ;
	double x_rho(eta_rho, xi_rho) ;
		x_rho:long_name = "x location of RHO-points" ;
		x_rho:units = "meter" ;
	double y_rho(eta_rho, xi_rho) ;
		y_rho:long_name = "y location of RHO-points" ;
		y_rho:units = "meter" ;
	double x_psi(eta_psi, xi_psi) ;
		x_psi:long_name = "x location of PSI-points" ;
		x_psi:units = "meter" ;
	double y_psi(eta_psi, xi_psi) ;
		y_psi:long_name = "y location of PSI-points" ;
		y_psi:units = "meter" ;
	double x_u(eta_u, xi_u) ;
		x_u:long_name = "x location of U-points" ;
		x_u:units = "meter" ;
	double y_u(eta_u, xi_u) ;
		y_u:long_name = "y location of U-points" ;
		y_u:units = "meter" ;
	double x_v(eta_v, xi_v) ;
		x_v:long_name = "x location of V-points" ;
		x_v:units = "meter" ;
	double y_v(eta_v, xi_v) ;
		y_v:long_name = "y location of V-points" ;
		y_v:units = "meter" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
	double lat_psi(eta_psi, xi_psi) ;
		lat_psi:long_name = "latitude of PSI-points" ;
		lat_psi:units = "degree_north" ;
	double lon_psi(eta_psi, xi_psi) ;
		lon_psi:long_name = "longitude of PSI-points" ;
		lon_psi:units = "degree_east" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:option\(0\) = "land" ;
		mask_rho:option\(1\) = "water" ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:option\(0\) = "land" ;
		mask_u:option\(1\) = "water" ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:option\(0\) = "land" ;
		mask_v:option\(1\) = "water" ;
	double mask_psi(eta_psi, xi_psi) ;
		mask_psi:long_name = "mask on PSI-points" ;
		mask_psi:option\(0\) = "land" ;
		mask_psi:option\(1\) = "water" ;
	double angle(eta_rho, xi_rho) ;
		angle:long_name = "angle between xi axis and east" ;
		angle:units = "radian" ;
	double N ;
		N:long_name = "Number of vertical layers" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
}
