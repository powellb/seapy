netcdf ini_hydro {

dimensions:
    xi_rho = 130 ;
    xi_u = 129 ;
    xi_v = 130 ;
    eta_rho = 130 ;
    eta_u = 130 ;
    eta_v = 129 ;
    s_rho = 20 ;
    s_w = 21 ;
    ocean_time = UNLIMITED ; // (0 currently)

variables:
  int Vtransform ;
    Vtransform:long_name = "vertical terrain-following transformation equation" ;
  int Vstretching ;
    Vstretching:long_name = "vertical terrain-following stretching function" ;
  double theta_s ;
    theta_s:long_name = "S-coordinate surface control parameter" ;
  double theta_b ;
    theta_b:long_name = "S-coordinate bottom control parameter" ;
  double Tcline ;
    Tcline:long_name = "S-coordinate surface/bottom layer width" ;
    Tcline:units = "meter" ;
  double hc ;
    hc:long_name = "S-coordinate parameter, critical depth" ;
    hc:units = "meter" ;
  double s_rho(s_rho) ;
    s_rho:long_name = "S-coordinate at RHO-points" ;
    s_rho:valid_min = -1. ;
    s_rho:valid_max = 0. ;
    s_rho:positive = "up" ;
    s_rho:standard_name = "ocean_s_coordinate_g1" ;
    s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
  double Cs_r(s_rho) ;
    Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
    Cs_r:valid_min = -1. ;
    Cs_r:valid_max = 0. ;
  double h(eta_rho, xi_rho) ;
    h:long_name = "bathymetry at RHO-points" ;
    h:units = "meter" ;
    h:coordinates = "lon_rho lat_rho" ;
  double angle(eta_rho, xi_rho) ;
      angle:long_name = "angle between xi axis and east" ;
      angle:units = "radian" ;
  double lon_rho(eta_rho, xi_rho) ;
    lon_rho:long_name = "longitude of RHO-points" ;
    lon_rho:units = "degree_east" ;
    lon_rho:standard_name = "longitude" ;
  double lat_rho(eta_rho, xi_rho) ;
    lat_rho:long_name = "latitude of RHO-points" ;
    lat_rho:units = "degree_north" ;
    lat_rho:standard_name = "latitude" ;
  double lon_u(eta_u, xi_u) ;
    lon_u:long_name = "longitude of U-points" ;
    lon_u:units = "degree_east" ;
    lon_u:standard_name = "longitude" ;
  double lat_u(eta_u, xi_u) ;
    lat_u:long_name = "latitude of U-points" ;
    lat_u:units = "degree_north" ;
    lat_u:standard_name = "latitude" ;
  double lon_v(eta_v, xi_v) ;
    lon_v:long_name = "longitude of V-points" ;
    lon_v:units = "degree_east" ;
    lon_v:standard_name = "longitude" ;
  double lat_v(eta_v, xi_v) ;
    lat_v:long_name = "latitude of V-points" ;
    lat_v:units = "degree_north" ;
    lat_v:standard_name = "latitude" ;
  double ocean_time(ocean_time) ;
      ocean_time:long_name = "time since initialization" ;
      ocean_time:units = "seconds since 0000-01-01 00:00:00" ;
  float zeta(ocean_time, eta_rho, xi_rho) ;
      zeta:long_name = "free-surface" ;
      zeta:units = "meter" ;
      zeta:coordinates = "lon_rho lat_rho ocean_time" ;
  float ubar(ocean_time, eta_u, xi_u) ;
      ubar:long_name = "vertically integrated u-momentum component" ;
      ubar:units = "meter second-1" ;
      ubar:coordinates = "lon_u lat_u ocean_time" ;
  float vbar(ocean_time, eta_v, xi_v) ;
      vbar:long_name = "vertically integrated v-momentum component" ;
      vbar:units = "meter second-1" ;
      vbar:coordinates = "lon_v lat_v ocean_time" ;
  float u(ocean_time, s_rho, eta_u, xi_u) ;
      u:long_name = "u-momentum component" ;
      u:units = "meter second-1" ;
      u:coordinates = "lon_u lat_u s_rho ocean_time" ;
  float v(ocean_time, s_rho, eta_v, xi_v) ;
      v:long_name = "v-momentum component" ;
      v:units = "meter second-1" ;
      v:coordinates = "lon_v lat_v s_rho ocean_time" ;
  float temp(ocean_time, s_rho, eta_rho, xi_rho) ;
      temp:long_name = "potential temperature" ;
      temp:units = "Celsius" ;
      temp:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float salt(ocean_time, s_rho, eta_rho, xi_rho) ;
      salt:long_name = "salinity" ;
      salt:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float alk(ocean_time, s_rho, eta_rho, xi_rho) ;
      alk:long_name = "Alkalinity" ;
      alk:units = "mol/kg" ;
      alk:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float cadet_arag(ocean_time, s_rho, eta_rho, xi_rho) ;
      cadet_arag:long_name = "Detrital Aragonite CaCO3" ;
      cadet_arag:units = "mol/kg" ;
      cadet_arag:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float cadet_calc(ocean_time, s_rho, eta_rho, xi_rho) ;
      cadet_calc:long_name = "Detrital Calcite CaCO3" ;
      cadet_calc:units = "mol/kg" ;
      cadet_calc:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float dic(ocean_time, s_rho, eta_rho, xi_rho) ;
      dic:long_name = "Dissolved Inorganic Carbon" ;
      dic:units = "mol/kg" ;
      dic:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float fed(ocean_time, s_rho, eta_rho, xi_rho) ;
      fed:long_name = "Dissolved Iron" ;
      fed:units = "mol/kg" ;
      fed:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float fedet(ocean_time, s_rho, eta_rho, xi_rho) ;
      fedet:long_name = "Detrital Iron" ;
      fedet:units = "mol/kg" ;
      fedet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float fedi(ocean_time, s_rho, eta_rho, xi_rho) ;
      fedi:long_name = "Diazotroph Iron" ;
      fedi:units = "mol/kg" ;
      fedi:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float felg(ocean_time, s_rho, eta_rho, xi_rho) ;
      felg:long_name = "Large Phytoplankton Iron" ;
      felg:units = "mol/kg" ;
      felg:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float fesm(ocean_time, s_rho, eta_rho, xi_rho) ;
      fesm:long_name = "Small Phytoplankton Iron" ;
      fesm:units = "mol/kg" ;
      fesm:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float ldon(ocean_time, s_rho, eta_rho, xi_rho) ;
      ldon:long_name = "Labile DON" ;
      ldon:units = "mol/kg" ;
      ldon:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float ldop(ocean_time, s_rho, eta_rho, xi_rho) ;
      ldop:long_name = "Labile DOP" ;
      ldop:units = "mol/kg" ;
      ldop:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float lith(ocean_time, s_rho, eta_rho, xi_rho) ;
      lith:long_name = "Lithogenic Aluminosilicate" ;
      lith:units = "g/kg" ;
      lith:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float lithdet(ocean_time, s_rho, eta_rho, xi_rho) ;
      lithdet:long_name = "Lithogenic Aluminosilicate, detrital" ;
      lithdet:units = "g/kg" ;
      lithdet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float nbact(ocean_time, s_rho, eta_rho, xi_rho) ;
      nbact:long_name = "Bacterial Nitrogen" ;
      nbact:units = "mol/kg" ;
      nbact:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float ndet(ocean_time, s_rho, eta_rho, xi_rho) ;
      ndet:long_name = "Detrital Nitrogen" ;
      ndet:units = "mol/kg" ;
      ndet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float ndi(ocean_time, s_rho, eta_rho, xi_rho) ;
      ndi:long_name = "Diazotroph Nitrogen" ;
      ndi:units = "mol/kg" ;
      ndi:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float nlg(ocean_time, s_rho, eta_rho, xi_rho) ;
      nlg:long_name = "Large Phytoplankton Nitrogen" ;
      nlg:units = "mol/kg" ;
      nlg:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float nsm(ocean_time, s_rho, eta_rho, xi_rho) ;
      nsm:long_name = "Small Phytoplankton Nitrogen" ;
      nsm:units = "mol/kg" ;
      nsm:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float nh4(ocean_time, s_rho, eta_rho, xi_rho) ;
      nh4:long_name = "Ammonia" ;
      nh4:units = "mol/kg" ;
      nh4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float no3(ocean_time, s_rho, eta_rho, xi_rho) ;
      no3:long_name = "Nitrate" ;
      no3:units = "mol/kg" ;
      no3:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float o2(ocean_time, s_rho, eta_rho, xi_rho) ;
      o2:long_name = "Oxygen" ;
      o2:units = "mol/kg" ;
      o2:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float pdet(ocean_time, s_rho, eta_rho, xi_rho) ;
      pdet:long_name = "Detrital Phosphorus" ;
      pdet:units = "mol/kg" ;
      pdet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float po4(ocean_time, s_rho, eta_rho, xi_rho) ;
      po4:long_name = "Phosphate" ;
      po4:units = "mol/kg" ;
      po4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float srdon(ocean_time, s_rho, eta_rho, xi_rho) ;
      srdon:long_name = "Semi-Refractory DON" ;
      srdon:units = "mol/kg" ;
      srdon:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float srdop(ocean_time, s_rho, eta_rho, xi_rho) ;
      srdop:long_name = "Semi-Refractory DOP" ;
      srdop:units = "mol/kg" ;
      srdop:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float sldon(ocean_time, s_rho, eta_rho, xi_rho) ;
      sldon:long_name = "Semilabile DON" ;
      sldon:units = "mol/kg" ;
      sldon:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float sldop(ocean_time, s_rho, eta_rho, xi_rho) ;
      sldop:long_name = "Semilabile DOP" ;
      sldop:units = "mol/kg" ;
      sldop:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float sidet(ocean_time, s_rho, eta_rho, xi_rho) ;
      sidet:long_name = "Detrital Silicon" ;
      sidet:units = "mol/kg" ;
      sidet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float silg(ocean_time, s_rho, eta_rho, xi_rho) ;
      silg:long_name = "Large Phytoplankton Silicon" ;
      silg:units = "mol/kg" ;
      silg:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float sio4(ocean_time, s_rho, eta_rho, xi_rho) ;
      sio4:long_name = "Silicate" ;
      sio4:units = "mol/kg" ;
      sio4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float nsmz(ocean_time, s_rho, eta_rho, xi_rho) ;
      nsmz:long_name = "Small Zooplankton Nitrogen" ;
      nsmz:units = "mol/kg" ;
      nsmz:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float nmdz(ocean_time, s_rho, eta_rho, xi_rho) ;
      nmdz:long_name = "Medium-sized Zooplankton Nitrogen" ;
      nmdz:units = "mol/kg" ;
      nmdz:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
  float nlgz(ocean_time, s_rho, eta_rho, xi_rho) ;
      nlgz:long_name = "Large Zooplankton Nitrogen" ;
      nlgz:units = "mol/kg" ;
      nlgz:coordinates = "lon_rho lat_rho s_rho ocean_time" ;

// global attributes:
        :type = "INITIALIZATION file" ;
}
