netcdf s4dvar_obs {

dimensions:
  survey = 1 ;
  state_variable = 20 ;
  datum = UNLIMITED ; // (0 currently)
variables:
  int spherical ;
    spherical:long_name = "grid type logical switch" ;
    spherical:flag_values = "0, 1" ;
    spherical:flag_meanings = "Cartesian spherical" ;
  int Nobs(survey) ;
    Nobs:long_name = "number of observations with the same survey time" ;
  double survey_time(survey) ;
    survey_time:long_name = "survey time" ;
    survey_time:units = "day" ;
  double obs_variance(state_variable) ;
    obs_variance:long_name = "global time and space observation variance" ;
    obs_variance:units = "squared state variable units" ;
  int obs_type(datum) ;
    obs_type:long_name = "model state variable associated with observation" ;
    obs_type:flag_values = "see global state variables" ;
  int obs_provenance(datum) ;
    obs_provenance:long_name = "observation origin" ;
  double obs_time(datum) ;
    obs_time:long_name = "time of observation" ;
    obs_time:units = "day" ;
  double obs_lat(datum) ;
    obs_lat:long_name = "latitude of observation" ;
    obs_lat:units = "degrees" ;
  double obs_lon(datum) ;
    obs_lon:long_name = "longitude of observation" ;
    obs_lon:units = "degrees" ;
  double obs_depth(datum) ;
    obs_depth:long_name = "depth of observation" ;
    obs_depth:units = "meter" ;
    obs_depth:negative = "downwards" ;
  double obs_Xgrid(datum) ;
    obs_Xgrid:long_name = "x-grid observation location" ;
    obs_Xgrid:left = "INT(obs_Xgrid(datum))" ;
    obs_Xgrid:right = "INT(obs_Xgrid(datum))+1" ;
  double obs_Ygrid(datum) ;
    obs_Ygrid:long_name = "y-grid observation location" ;
    obs_Ygrid:top = "INT(obs_Ygrid(datum))+1" ;
    obs_Ygrid:bottom = "INT(obs_Ygrid(datum))" ;
  double obs_Zgrid(datum) ;
    obs_Zgrid:long_name = "z-grid observation location" ;
    obs_Zgrid:up = "INT(obs_Zgrid(datum))+1" ;
    obs_Zgrid:down = "INT(obs_Zgrid(datum))" ;
  double obs_error(datum) ;
    obs_error:long_name = "observation error covariance" ;
    obs_error:units = "squared state variable units" ;
  double obs_value(datum) ;
    obs_value:long_name = "observation value" ;
    obs_value:units = "state variable units" ;
  double obs_meta(datum) ;
    obs_meta:long_name = "observation meta value" ;
    obs_meta:units = "observational secondary units" ;

// global attributes:
    :type = "ROMS Observations" ;
}
